module line_drawing_FSM (clk, start);
	input clk, start, 
	

	 
endmodule 