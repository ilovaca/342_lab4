module line_drawing_datapath ();

	register_nbit #(.SIZE(9)) x0 ();
	register_nbit #(.SIZE(9)) x1 ();
	register_nbit #(.SIZE(8)) y0 ();
	register_nbit #(.SIZE(8)) y1 ();
	register_nbit #(.SIZE(9)) 
endmodule